library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity project_reti_logiche is
    port(
        i_clk       : in std_logic;
        i_rst       : in std_logic;
        i_start     : in std_logic;
        i_data      : in std_logic_vector(7 downto 0);
        o_address   : out std_logic_vector(15 downto 0);
        o_done      : out std_logic;
        o_en        : out std_logic;
        o_we        : out std_logic;
        o_data      : out std_logic_vector(7 downto 0)
    );
end project_reti_logiche;

architecture rtl of project_reti_logiche is
    signal N_COL, N_RIG : unsigned(7 downto 0);
    signal COUNTER, J : unsigned(15 downto 0);
    signal DELTA_VALUE, MAX_PIXEL_VALUE, MIN_PIXEL_VALUE, TEMP_PIXEL, NEW_PIXEL_VALUE, CURRENT_PIXEL_VALUE, BEFORE_SHIFT : unsigned(7 downto 0);
    signal TOT_PIXEL, K , TOT_PIXEL_ORIGINAL: unsigned(15 downto 0);
    signal SHIFT_LEVEL: integer;
    signal OverFlow, IsClean, synced : std_logic := '0';

    type t_state is (FIRST, RESET, WAITING, START, READCOL, READRIG, LOADTOT, MAXMIN, LOADDELTA, LOADSHIFT, CALCULATENEWVALUE, HASOVERFLOWED, WRITENEWVALUE, SYNC, DONE);
    signal state : t_state;
    
    begin
        process(i_clk)
        begin
            if rising_edge(i_clk) then
                if i_rst = '1'  and isClean = '0' then
                    state <= RESET;
                end if;
            
                if state = RESET then
                    if synced = '0' then
                        synced <= '1';
                    else
                        if IsClean = '0' then
                            N_COL <= (others => '0');
                            N_RIG <= (others => '0');
                            DELTA_VALUE <= (others => '0');
                            MAX_PIXEL_VALUE <= (others => '0');
                            MIN_PIXEL_VALUE <= (others => '1');
                            TEMP_PIXEL <= (others => '0');
                            NEW_PIXEL_VALUE <= (others => '0');
                            CURRENT_PIXEL_VALUE <= (others => '0');
                            COUNTER <= (others => '0');
                            J <= (others => '0');
                            TOT_PIXEL_ORIGINAL <= (others => '0');
                            TOT_PIXEL <= (others => '0');
                            SHIFT_LEVEL <= 0;
                            K <= (others => '0');
                            TOT_PIXEL <= (others => '0');
                            BEFORE_SHIFT <= "00000000";
                            o_en <= '0';
                            o_we <= '0';
                            o_done <= '0';
                            o_address <= (others => '0');
                            o_data <= (others => '0');
                            OverFlow <= '0';
                            synced <= '0';
                            IsClean <= '1';
                            report "initialized";
                            
                            state <= WAITING;
                        end if;
                    end if;
                
                elsif state = WAITING then
                    if synced = '0' then
                        synced <= '1';
                    elsif i_start = '1' then
                        state <= START;
                        o_en <= '1';
                        synced <= '0';
                    end if;
                
                elsif state = START then
                    if synced = '0' then
                        synced <= '1';
                    else
                        state <= READCOL;
                        o_address <= std_logic_vector(COUNTER);
                        COUNTER <= J + 1;
                        J <= COUNTER + 1;
                        isClean <= '0';
                        synced <= '0';
                    end if;
                
                elsif state = READCOL then
                    if synced = '0' then
                        synced <= '1';
                    else
                        N_COL <= unsigned(i_data);
                        state <= READRIG;
                        
                        o_address <= std_logic_vector(COUNTER);
                        COUNTER <= J + 1;
                        J <= COUNTER + 1;
                        
                        synced <= '0';
                    end if;
                
                
                elsif state = READRIG then
                    if synced = '0' then
                        synced <= '1';
                    else
                        N_RIG <= unsigned(i_data);
                        state <= LOADTOT;
                        synced <= '0';
                    end if;
                
                elsif state = LOADTOT then
                    if synced = '0' then
                        synced <= '1';
                    else
                        TOT_PIXEL <= (N_COL * N_RIG);
                        TOT_PIXEL_ORIGINAL <= (N_COL * N_RIG);
                        K <= (N_COL * N_RIG);
                        
                        o_address <= std_logic_vector(COUNTER);
                        COUNTER <= J + 1;
                        J <= COUNTER + 1;
                        
                        state <= MAXMIN;
                        synced <= '0';
                    end if;
                
                elsif state = MAXMIN then
                    if synced = '0' then
                        synced <= '1';
                    else
                        if TOT_PIXEL > 0 then
                            CURRENT_PIXEL_VALUE  <= unsigned(i_data);--ce lo possiamo risparmiare, � per vedere meglio la simulazione
                            if unsigned(i_data) > MAX_PIXEL_VALUE then
                                MAX_PIXEL_VALUE  <= unsigned(i_data);
                            end if; 
                            
                            if unsigned(i_data) < MIN_PIXEL_VALUE then
                                MIN_PIXEL_VALUE  <= unsigned(i_data);
                            end if;
                            
                            o_address <= std_logic_vector(COUNTER);
                            COUNTER <= J + 1;
                            J <= COUNTER + 1;
                           
                            TOT_PIXEL <= K - 1;
                            K <= TOT_PIXEL - 1;
                        else 
                            state <= LOADDELTA;
                        end if;
                        synced <= '0';
                    end if;
                
                elsif state = LOADDELTA then
                    if synced = '0' then
                        synced <= '1';
                    else
                        DELTA_VALUE <= MAX_PIXEL_VALUE - MIN_PIXEL_VALUE;
                        COUNTER <= (others => '0');
                        COUNTER(1) <= '1';
                        J <= (others => '0');
                        J(1) <= '1';
                        state <= LOADSHIFT;
                        synced <= '0';
                    end if;
                
                elsif state = LOADSHIFT then
                if synced = '0' then
                        synced <= '1';
                    else
                        TOT_PIXEL <= TOT_PIXEL_ORIGINAL;
                        K <= TOT_PIXEL_ORIGINAL;
                        if DELTA_VALUE = "00000000" then
                            SHIFT_LEVEL <= 8;
                        elsif  (DELTA_VALUE="00000001" or DELTA_VALUE="00000010") then
                            SHIFT_LEVEL <= 7;
                        elsif  (DELTA_VALUE>="00000011" and DELTA_VALUE<="00000110") then
                            SHIFT_LEVEL <= 6;
                        elsif  (DELTA_VALUE>="00000111" and DELTA_VALUE<="00001110") then
                            SHIFT_LEVEL <= 5;
                        elsif  (DELTA_VALUE>="00001111" and DELTA_VALUE<="00011110") then
                            SHIFT_LEVEL <= 4;                                                                        
                        elsif  (DELTA_VALUE>="00011111" and DELTA_VALUE<="00111110") then
                            SHIFT_LEVEL <= 3;
                        elsif  (DELTA_VALUE>="00111111" and DELTA_VALUE<="01111110") then
                            SHIFT_LEVEL <= 2;
                        elsif  (DELTA_VALUE>="01111111" and DELTA_VALUE<="11111110") then
                            SHIFT_LEVEL <= 1;  
                        elsif  DELTA_VALUE="11111111" then
                            SHIFT_LEVEL <= 0;                                                               
                        end if;
                        
                        state <= CALCULATENEWVALUE;
                        o_address <= std_logic_vector(COUNTER);
                        synced <= '0';
                    end if;
                
                elsif state = CALCULATENEWVALUE then
                    if synced = '0' then
                        synced <= '1';
                    else
                        if TOT_PIXEL > 0 then
                            BEFORE_SHIFT <= unsigned(i_data) - MIN_PIXEL_VALUE;
                            TEMP_PIXEL <= shift_left((unsigned(i_data) - MIN_PIXEL_VALUE), SHIFT_LEVEL);
                            TOT_PIXEL <= K - 1;
                            K <= TOT_PIXEL - 1;
                            
                            o_address <= std_logic_vector(COUNTER + TOT_PIXEL_ORIGINAL );
                            COUNTER <= J + 1;
                            J <= COUNTER + 1;
                            
                            state <= HASOVERFLOWED;
                        else 
                            state <= DONE;
                        end if;
                        synced <= '0';
                    end if;
                
                elsif state = HASOVERFLOWED then
                    if synced = '0' then
                        synced <= '1';
                    else
                        if SHIFT_LEVEL > 0 then
                            if(SHIFT_LEVEL = 7) then
                                for i in 7 downto 1 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            elsif(SHIFT_LEVEL = 6) then
                                for i in 7 downto 2 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            elsif(SHIFT_LEVEL = 5) then
                                for i in 7 downto 3 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            elsif(SHIFT_LEVEL = 4) then
                                for i in 7 downto 4 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            elsif(SHIFT_LEVEL = 3) then
                                for i in 7 downto 5 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            elsif(SHIFT_LEVEL = 2) then
                                for i in 7 downto 6 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            elsif(SHIFT_LEVEL = 1) then
                                for i in 7 downto 7 loop
                                    if(BEFORE_SHIFT(i) = '1' and OverFlow = '0') then
                                        OverFlow <= '1';
                                    end if;
                                end loop;
                            end if;
                        end if;
                        state <= WRITENEWVALUE;
                        o_we <= '1';
                        synced <= '0';
                    end if;
                
                elsif state = WRITENEWVALUE then
                    if synced = '0' then
                        synced <= '1';
                    else
                        if OverFlow = '1' then
                            o_data <= "11111111";
                        else
                            o_data <= std_logic_vector(TEMP_PIXEL);
                        end if;
                        OverFlow <= '0';
                        state <= SYNC;
                        synced <= '0';
                    end if;
                    
                elsif state = SYNC then
                    if synced = '0' then
                        synced <= '1';
                    else
                        state <= CALCULATENEWVALUE;
                        o_address <= std_logic_vector(COUNTER);
                        o_we <= '0';
                        synced <= '0';
                    end if;
                
                elsif state = DONE then
                    if synced = '0' then
                        synced <= '1';
                    else
                        if i_start = '1' then
                            o_done <= '1';
                            o_en <= '0';
                        elsif i_start = '0' then
                            o_done <= '0';
                            state <= RESET;
                        end if;
                        synced <= '0';
                    end if;
                
                end if;
            end if;
        end process;
end architecture;